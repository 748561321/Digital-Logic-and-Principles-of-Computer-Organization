module bcd7seg(
	input [7:0] b,
	output reg [6:0] h1,
	output reg [6:0] h2
);

	always @(b) begin
		if(b==8'h00)begin
			h1=7'b1111111;
			h2=7'b1111111;
		end
		else begin
			case(b[3:0])
			4'b0000:h1=7'b1000000;
			4'b0001:h1=7'b1111001;
			4'b0010:h1=7'b0100100;
			4'b0011:h1=7'b0110000;
			4'b0100:h1=7'b0011001;
			4'b0101:h1=7'b0010010;
			4'b0110:h1=7'b0000010;
			4'b0111:h1=7'b1111000;
			4'b1000:h1=7'b0000000;
			4'b1001:h1=7'b0011000;
			4'b1010:h1=7'b0001000;
			4'b1011:h1=7'b0000011;
			4'b1100:h1=7'b1000110;
			4'b1101:h1=7'b0100001;
			4'b1110:h1=7'b0000110;
			4'b1111:h1=7'b0001110;
			endcase
			casex(b[7:4])
			4'b0000:h2=7'b1000000;
			4'b0001:h2=7'b1111001;
			4'b0010:h2=7'b0100100;
			4'b0011:h2=7'b0110000;
			4'b0100:h2=7'b0011001;
			4'b0101:h2=7'b0010010;
			4'b0110:h2=7'b0000010;
			4'b0111:h2=7'b1111000;
			4'b1000:h2=7'b0000000;
			4'b1001:h2=7'b0011000;
			4'b1010:h2=7'b0001000;
			4'b1011:h2=7'b0000011;
			4'b1100:h2=7'b1000110;
			4'b1101:h2=7'b0100001;
			4'b1110:h2=7'b0000110;
			4'b1111:h2=7'b0001110;
			endcase
		end
	end

endmodule